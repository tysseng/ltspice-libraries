POT1.CIR - POTENTIOMETER
*
* WIPER POSITION: 0V=CCW, 1V=CW
VPOS	20	0	PWL(0MS 0V   100MS 1V)
RPOS	20	0	1MEG
*
* OFFSET VOLTAGE TRIM
VS	10	0	10V
R1	10	11	9K
XPOT1	0 12 11	20 0	POT_1K
RL	12	0	100K
*
* RESISTANCE VALUE TRIM
IS	0	15	1A
XPOT2	15 16	16 20 0 POT_1K
R2	16	0	19.5K
*
*
* POTENTIOMETER SUBCIRCUIT
*
* TERMINALS:	1-CCW , 2-WIPER, 3-CW 
* WIPER POSITION VOLTAGE:	7-POS,8-NEG
*
.SUBCKT POT_1K   1 2 3  7 8 
E_RA	1 4	 VALUE = { V(7,8) * 1K * I(VSENSE1) }
VSENSE1	4	5	DC	0V
RS	5	2	1
E_RB	5 6	 VALUE = { (1-V(7,8)) * 1K * I(VSENSE2) }
VSENSE2	6	3	DC	0V
.ENDS
*
*
* ANALYSIS
.TRAN 	0.1MS  100MS
* VIEW RESULTS
.PRINT	TRAN 	V(12)
.PROBE
.END